* C:\Users\user\Documents\bjtinverters.sch

* Schematics Version 9.1 - Web Update 1
* Thu Jul 12 00:00:05 2018



** Analysis setup **
.DC LIN V_Vin 0 100 1 
.MC 50 DC V([Vout]) YMAX
+  OUTPUT ALL
.OP 
.LIB "C:\Users\user\Documents\bjtinverters.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "bjtinverters.net"
.INC "bjtinverters.als"


.probe


.END
